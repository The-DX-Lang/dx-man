module string_parser

pub fn identity_parser(input string) ?string {
	return input
}
